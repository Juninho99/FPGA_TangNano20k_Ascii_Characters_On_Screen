//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sun Sep 24 16:22:42 2023

module Gowin_pROM_ascii (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h000000007E818199BD8181A5817E000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000010387CFEFEFEFE6C00000000000000007EFFFFE7C3FFFFDBFF7E0000;
defparam prom_inst_0.INIT_RAM_02 = 256'h000000003C1818E7E7E73C3C18000000000000000010387CFE7C381000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000000000183C3C18000000000000000000003C18187EFFFF7E3C18000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h00000000003C664242663C0000000000FFFFFFFFFFFFE7C3C3E7FFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000078CCCCCCCC78321A0E1E0000FFFFFFFFFFC399BDBD99C3FFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'h00000000E0F070303030303F333F00000000000018187E183C666666663C0000;
defparam prom_inst_0.INIT_RAM_07 = 256'h000000001818DB3CE73CDB1818000000000000C0E6E767636363637F637F0000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000002060E1E3EFE3E1E0E0602000000000080C0E0F0F8FEF8F0E0C08000;
defparam prom_inst_0.INIT_RAM_09 = 256'h000000006666006666666666666600000000000000183C7E1818187E3C180000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000007CC60C386CC6C66C3860C67C00000000001B1B1B1B1B7BDBDBDB7F0000;
defparam prom_inst_0.INIT_RAM_0B = 256'h000000307E183C7E1818187E3C18000000000000FEFEFEFE0000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h00000000183C7E18181818181818000000000000181818181818187E3C180000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000003060FE60300000000000000000000000180CFE0C180000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000002466FF66240000000000000000000000FEC0C0C0000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000001038387C7CFEFE000000000000000000FEFE7C7C38381000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h000000001818001818183C3C3C18000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h000000006C6CFE6C6C6CFE6C6C00000000000000000000000000002466666600;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000086C66030180CC6C200000000000018187CC68606067CC0C2C67C1818;
defparam prom_inst_0.INIT_RAM_13 = 256'h000000000000000000000060303030000000000076CCCCCCDC76386C6C380000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000030180C0C0C0C0C0C18300000000000000C18303030303030180C0000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000000018187E18180000000000000000000000663CFF3C660000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000000000007E0000000000000000000030181818000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000080C06030180C06020000000000000000181800000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h000000007E1818181818187838180000000000007CC6C6E6F6DECEC6C67C0000;
defparam prom_inst_0.INIT_RAM_19 = 256'h000000007CC60606063C0606C67C000000000000FEC6C06030180C06C67C0000;
defparam prom_inst_0.INIT_RAM_1A = 256'h000000007CC6060606FCC0C0C0FE0000000000001E0C0C0CFECC6C3C1C0C0000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000030303030180C0606C6FE0000000000007CC6C6C6C6FCC0C060380000;
defparam prom_inst_0.INIT_RAM_1C = 256'h00000000780C0606067EC6C6C67C0000000000007CC6C6C6C67CC6C6C67C0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000030181800000018180000000000000000001818000000181800000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h000000000000007E00007E000000000000000000060C18306030180C06000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h000000001818001818180CC6C67C0000000000006030180C060C183060000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h00000000C6C6C6C6FEC6C66C38100000000000007CC0DCDEDEDEC6C6C67C0000;
defparam prom_inst_0.INIT_RAM_21 = 256'h000000003C66C2C0C0C0C0C2663C000000000000FC666666667C666666FC0000;
defparam prom_inst_0.INIT_RAM_22 = 256'h00000000FE6662606878686266FE000000000000F86C6666666666666CF80000;
defparam prom_inst_0.INIT_RAM_23 = 256'h000000003A66C6C6DEC0C0C2663C000000000000F06060606878686266FE0000;
defparam prom_inst_0.INIT_RAM_24 = 256'h000000003C18181818181818183C000000000000C6C6C6C6C6FEC6C6C6C60000;
defparam prom_inst_0.INIT_RAM_25 = 256'h00000000E666666C78786C6666E600000000000078CCCCCC0C0C0C0C0C1E0000;
defparam prom_inst_0.INIT_RAM_26 = 256'h00000000C3C3C3C3C3DBFFFFE7C3000000000000FE6662606060606060F00000;
defparam prom_inst_0.INIT_RAM_27 = 256'h000000007CC6C6C6C6C6C6C6C67C000000000000C6C6C6C6CEDEFEF6E6C60000;
defparam prom_inst_0.INIT_RAM_28 = 256'h00000E0C7CDED6C6C6C6C6C6C67C000000000000F0606060607C666666FC0000;
defparam prom_inst_0.INIT_RAM_29 = 256'h000000007CC6C6060C3860C6C67C000000000000E66666666C7C666666FC0000;
defparam prom_inst_0.INIT_RAM_2A = 256'h000000007CC6C6C6C6C6C6C6C6C60000000000003C18181818181899DBFF0000;
defparam prom_inst_0.INIT_RAM_2B = 256'h000000006666FFDBDBC3C3C3C3C3000000000000183C66C3C3C3C3C3C3C30000;
defparam prom_inst_0.INIT_RAM_2C = 256'h000000003C181818183C66C3C3C3000000000000C3C3663C18183C66C3C30000;
defparam prom_inst_0.INIT_RAM_2D = 256'h000000003C30303030303030303C000000000000FFC3C16030180C86C3FF0000;
defparam prom_inst_0.INIT_RAM_2E = 256'h000000003C0C0C0C0C0C0C0C0C3C00000000000002060E1C3870E0C080000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000FF00000000000000000000000000000000000000000000000000C66C3810;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000076CCCCCC7C0C78000000000000000000000000000000000000183030;
defparam prom_inst_0.INIT_RAM_31 = 256'h000000007CC6C0C0C0C67C0000000000000000007C666666666C786060E00000;
defparam prom_inst_0.INIT_RAM_32 = 256'h000000007CC6C0C0FEC67C00000000000000000076CCCCCCCC6C3C0C0C1C0000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0078CC0C7CCCCCCCCCCC76000000000000000000F060606060F060646C380000;
defparam prom_inst_0.INIT_RAM_34 = 256'h000000003C181818181838001818000000000000E666666666766C6060E00000;
defparam prom_inst_0.INIT_RAM_35 = 256'h00000000E6666C78786C666060E00000003C66660606060606060E0006060000;
defparam prom_inst_0.INIT_RAM_36 = 256'h00000000DBDBDBDBDBFFE60000000000000000003C1818181818181818380000;
defparam prom_inst_0.INIT_RAM_37 = 256'h000000007CC6C6C6C6C67C000000000000000000666666666666DC0000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h001E0C0C7CCCCCCCCCCC76000000000000F060607C6666666666DC0000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h000000007CC60C3860C67C000000000000000000F06060606676DC0000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000076CCCCCCCCCCCC0000000000000000001C3630303030FC3030100000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000066FFDBDBC3C3C3000000000000000000183C66C3C3C3C30000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h00F80C067EC6C6C6C6C6C6000000000000000000C3663C183C66C30000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h000000000E18181818701818180E000000000000FEC6603018CCFE0000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000070181818180E18181870000000000000181818181800181818180000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000FEC6C6C66C381000000000000000000000000000000000DC760000;

endmodule //Gowin_pROM_ascii
